library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package eth_pack is
    constant MAX_ETH_FRAME_SIZE : natural := 1530;
end package eth_pack;

package body eth_pack is

end package body eth_pack;